library ieee;
use ieee.std_logic_1164.all;

use ieee.numeric_std.all;

package pkg is
  type registers is array(natural range <>) of std_logic_vector(31 downto 0);
end package;

package body pkg is
end package body;