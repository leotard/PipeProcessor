library ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;



ENTITY HazardDetection IS
	port(
		flag : in std_logic;
		instruction: in std_logic_vector(31 downto 0);
		previous_inst: in std_logic_vector(31 downto 0);
		current_data_stall: in std_logic_vector(2 downto 0);
		stall: out std_logic_vector(2 downto 0)
	);
		
END HazardDetection;



ARCHITECTURE arch OF HazardDetection IS

--signal holds register number and number of stalls left (first 3 bits)
signal dest_reg_1, dest_reg_2, dest_reg_3, dest_reg_4, past_reg_1, past_reg_2: std_logic_vector(7 downto 0):="00011110";
signal past_stall : std_logic_vector(2 downto 0):="000";
signal temp : std_logic_vector(2 downto 0):="000";

constant R_TYPE : std_logic_vector(5 downto 0):= "000000";
constant ADDI : std_logic_vector(5 downto 0):= "001000";
constant slti : std_logic_vector(5 downto 0):= "001010";
constant LW : std_logic_vector(5 downto 0):= "100011";
constant BEQ : std_logic_vector(5 downto 0):= "000100";
constant BNE : std_logic_vector(5 downto 0):= "000101";


begin

process(instruction)


variable op_code : std_logic_vector(5 downto 0);
variable arg1, arg2, arg3: std_logic_vector(4 downto 0);
variable var_stall, var_past_stall: std_logic_vector(2 downto 0);
variable var_stall_temp_1, var_stall_temp_2 : std_logic_vector(2 downto 0);
variable var_dest_reg_1, var_dest_reg_2, var_dest_reg_3:std_logic_vector(7 downto 0);

begin

	op_code := instruction(31 downto 26);
	arg1 := instruction(25 downto 21);
	arg2 := instruction(20 downto 16);
	arg3 := instruction(15 downto 11);
	var_past_stall := std_logic_vector(to_unsigned(to_integer(unsigned(past_stall)) - 1, var_past_stall'length));
	if(instruction /= "00000000000000000000000000000000" AND previous_inst /= "00000000000000000000000000000000") then
			if(op_code = R_TYPE OR op_code = BNE OR op_code = BEQ) then
				if(arg3 /= "00000") then
					if(arg1 = dest_reg_1(4 downto 0)) then
						var_stall_temp_1 := dest_reg_1(7 downto 5);
					elsif(arg1 = dest_reg_2(4 downto 0)) then
						var_stall_temp_1 := dest_reg_2(7 downto 5);
					elsif(arg1 = dest_reg_3(4 downto 0)) then
						var_stall_temp_1 := dest_reg_3(7 downto 5);
					else 
						var_stall_temp_1 := "000";
					end if;
					if(arg2 = dest_reg_1(4 downto 0)) then
						var_stall_temp_2 := dest_reg_1(7 downto 5);
					elsif(arg2 = dest_reg_2(4 downto 0)) then
						var_stall_temp_2 := dest_reg_2(7 downto 5);
					elsif(arg2 = dest_reg_3(4 downto 0)) then
						var_stall_temp_2 := dest_reg_3(7 downto 5);
					else 
						var_stall_temp_2 := "000";
					end if;
					if(to_integer(unsigned(var_stall_temp_1)) > to_integer(unsigned(var_stall_temp_2))) then
						var_stall := var_stall_temp_1;
					else
						var_stall := var_stall_temp_2;
					end if;
					
					
				else
					if(past_stall /= "000") then
						var_stall := current_data_stall;
					else
						var_stall := "000";
					end if;
					
				end if;
			elsif(op_code = ADDI OR op_code = SLTI OR op_code = LW) then
				if(arg2 /= "00000") then
					if(arg1 = dest_reg_1(4 downto 0)) then
						var_stall_temp_1 := dest_reg_1(7 downto 5);
					elsif(arg1 = dest_reg_2(4 downto 0)) then
						var_stall_temp_1 := dest_reg_2(7 downto 5);
					elsif(arg1 = dest_reg_3(4 downto 0)) then
						var_stall_temp_1 := dest_reg_3(7 downto 5);
					else 
						var_stall_temp_1 := "000";
					end if;
					var_stall := var_stall_temp_1;
					
				else
					if(past_stall /= "000") then
						var_stall := current_data_stall;
					else
						var_stall := "000";
					end if;
					
				end if;
				--stall <= var_stall;
			end if;
	else
		if(past_stall /= "000") then
			var_stall := current_data_stall;
		else
			var_stall := "000";
		end if;
		
	end if;

	if(current_data_stall /= "000") then
		stall <= current_data_stall;
		past_stall <= current_data_stall;
	else
		stall <= var_stall;
		past_stall <= var_stall;
	end if;

	var_dest_reg_1 := dest_reg_1;
	var_dest_reg_2 := dest_reg_2;
	var_dest_reg_3 := dest_reg_3;
	dest_reg_2(4 downto 0) <= dest_reg_1(4 downto 0);
	dest_reg_3(4 downto 0) <= dest_reg_2(4 downto 0);
	if(dest_reg_1(7 downto 5) /= "000") then
		dest_reg_2(7 downto 5) <= std_logic_vector(to_unsigned(to_integer(unsigned(var_dest_reg_1(7 downto 5))) - 1, 3));
	end if;
	if(dest_reg_2(7 downto 5) /= "000") then
		dest_reg_3(7 downto 5) <= std_logic_vector(to_unsigned(to_integer(unsigned(var_dest_reg_2(7 downto 5))) - 1, 3));
	end if;
	
	if(instruction(31 downto 26) = R_TYPE AND instruction /= "00000000000000000000000000000000" AND instruction(5 downto 0) /="001000") then
		dest_reg_1(7 downto 5) <= "011";
		dest_reg_1(4 downto 0) <= instruction(15 downto 11);
	elsif(instruction(31 downto 26) = SLTI OR instruction(31 downto 26) = ADDI OR instruction(31 downto 26) = LW) then
		dest_reg_1(7 downto 5) <= "011";
		dest_reg_1(4 downto 0) <= instruction(20 downto 16);
	else
		dest_reg_1(4 downto 0) <= var_dest_reg_2(4 downto 0);
		dest_reg_2(4 downto 0) <= var_dest_reg_3(4 downto 0);
		--dest_reg_1 <= "00011111"; -- Store impossible register
	end if;

end process;
end arch;